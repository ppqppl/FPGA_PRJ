module PWM_Beep (
    output      wire        beep
);
    assign beep = 1'b0;
endmodule //beep