library verilog;
use verilog.vl_types.all;
entity pwn_tb is
end pwn_tb;
