module led (
    
);

endmodule //led