module KLED(
  input clk,
  input [3:0] key,
  output [3:0] led
);

  parameter MAX_COUNT = 26'd5000_0000; // 设定计数器的最大值

  reg [4:0] count_0, count_1, count_2, count_3; // 计数器
  reg [1:0] state_0, state_1, state_2, state_3; // 当前状态
  reg db_0, db_1, db_2, db_3; // 按键去抖动信号

  always @(posedge clk) begin
    if (key[0] != db_0) begin
      count_0 <= 0;
      db_0 <= key[0];
    end else if (count_0 == MAX_COUNT) begin
      db_0 <= key[0];
      if (db_0 == 1'b0) begin
        case (state_0)
          2'b00: state_0 <= 2'b01;
          2'b01: state_0 <= 2'b10;
          2'b10: state_0 <= 2'b11;
          2'b11: state_0 <= 2'b00;
        endcase
      end
    end else begin
      count_0 <= count_0 + 1;
    end

    if (key[1] != db_1) begin
      count_1 <= 0;
      db_1 <= key[1];
    end else if (count_1 == MAX_COUNT) begin
      db_1 <= key[1];
      if (db_1 == 1'b0) begin
        case (state_1)
          2'b00: state_1 <= 2'b01;
          2'b01: state_1 <= 2'b10;
          2'b10: state_1 <= 2'b11;
          2'b11: state_1 <= 2'b00;
        endcase
      end
    end else begin
      count_1 <= count_1 + 1;
    end

    if (key[2] != db_2) begin
      count_2 <= 0;
      db_2 <= key[2];
    end else if (count_2 == MAX_COUNT) begin
      db_2 <= key[2];
      if (db_2 == 1'b0) begin
        case (state_2)
          2'b00: state_2 <= 2'b01;
          2'b01: state_2 <= 2'b10;
          2'b10: state_2 <= 2'b11;
          2'b11: state_2 <= 2'b00;
        endcase
      end
    end else begin
      count_2 <= count_2 + 1;
    end

    if (key[3] != db_3) begin
      count_3 <= 0;
      db_3 <= key[3];
    end else if (count_3 == MAX_COUNT) begin
      db_3 <= key[3];
      if (db_3 == 1'b0) begin
        case (state_3)
          2'b00: state_3 <= 2'b01;
          2'b01: state_3 <= 2'b10;
          2'b10: state_3 <= 2'b11;
          2'b11: state_3 <= 2'b00;
        endcase
      end
    end else begin
      count_3 <= count_3 + 1;
    end
  end

  assign led[0] = (state_0[0] ^ state_0[1]);
  assign led[1] = (state_1[0] ^ state_1[1]);
  assign led[2] = (state_2[0] ^ state_2[1]);
  assign led[3] = (state_3[0] ^ state_3[1]);

endmodule