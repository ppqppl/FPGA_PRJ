module beep (
    
);

endmodule //beep