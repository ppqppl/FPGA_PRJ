module i2c_ctrl (
    input   wire    clk,
    input   wire    rst_n,

    output  wire    scl,
    inout   wire    sda 
);



endmodule //i2c_ctrl