module key (
    input   wire            clk     ,
    input   wire            rstn    ,
    input   wire    [3:0]   key_in  

);

endmodule //key